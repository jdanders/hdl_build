package pkg1;
  localparam PKG1 = 0;
endpackage: pkg1
