module submod2 (
  input wire bit_in,
  output wire bit_out
  );

  assign bit_out = bit_in;

endmodule: submod2
