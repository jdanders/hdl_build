package pkg2;
  localparam PKG2 = 0;
  function logic [1:0]  data_to_pipe (input data);
    return '0;
  endfunction: data_to_pipe

endpackage: pkg2
