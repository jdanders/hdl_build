localparam VALUE=1;
