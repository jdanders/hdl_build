package pkg2;
  localparam PKG2 = 0;
endpackage: pkg2
